
module file_reader_tb (  );
  wire   clk;

  CLKINVX8 U1 ( .A(clk), .Y(clk) );
endmodule

